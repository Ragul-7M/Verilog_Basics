module or_gate(
    input A,
    input B,
    output Y
    );
    or(Y,A,B);
endmodule
